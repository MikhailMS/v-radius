module protocol

